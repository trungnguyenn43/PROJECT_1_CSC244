
module NextStateLogic(
		input logic [3:0] S,
		input logic [1:0] A,
		
		output logic [3:0] Out
);
	
	logic [8:0] S_next;
	
	//Get next state
	assign S_next[0] = ~S[3] & ~S[2] & ~S[1] & ~S[0] & ~A[1] & ~A[0] //S0 -- 00
							| ~S[3] & S[2] & ~S[1] & S[0] & ~A[1] & ~A[0]  //S5 -- 00
							| ~S[3] & S[2] & S[1] & ~S[0] & ~A[1] & ~A[0]  //S6 -- 00
							| ~S[3] & S[2] & S[1] & S[0] & ~A[1] & ~A[0]  //S7 -- 00
							| S[3] & ~S[2] & ~S[1] & ~S[0] & ~A[1] & ~A[0]; //S8 -- 00
	
	assign S_next[1] = ~S[3] & ~S[2] & ~S[1] & ~S[0] & ~A[1] & A[0] //S0 - 01
							| ~S[3] & ~S[2] & ~S[1] & S[0] & ~A[1] & ~A[0] //S1 -- 00
							| ~S[3] & S[2] & ~S[1] & S[0] & ~A[1] & A[0]; //S5 - 01
	
	assign S_next[2] = ~S[3] & ~S[2] & ~S[1] & ~S[0] & A[1] & ~A[0] //S0 - 10
							| ~S[3] & ~S[2] & ~S[1] & S[0] & ~A[1] & A[0] //S1 -- 01
							| ~S[3] & ~S[2] & S[1] & ~S[0] & ~A[1] & ~A[0] //S2 - 00
							| ~S[3] & S[2] & S[1] & ~S[0] & ~A[1] & A[0]  //S6 -- 01
							| ~S[3] & S[2] & ~S[1] & S[0] & A[1] & ~A[0];  //S5 -- 10
							
	assign S_next[3] = ~S[3] & ~S[2] & ~S[1] & S[0] & A[1] & ~A[0] //S1 -- 10
							| ~S[3] & ~S[2] & S[1] & S[0] & ~A[1] & ~A[0] //S3 -- 00
							| ~S[3] & ~S[2] & S[1] & ~S[0] & ~A[1] & A[0] //S2 -- 01
							| ~S[3] & S[2] & S[1] & ~S[0] & A[1] & ~A[0] //S6 -- 10
							| ~S[3] & S[2] & S[1] & S[0] & ~A[1] & A[0]; //S7 -- 01
							
	assign S_next[4] = ~S[3] & ~S[2] & ~S[1] & ~S[0] & A[1] & A[0] //S0 -- 11
							| ~S[3] & ~S[2] & S[1] & S[0] & ~A[1] & A[0] //S3 -- 01
							| ~S[3] & ~S[2] & S[1] & ~S[0] & A[1] & ~A[0] //S2  -- 10
							| ~S[3] & S[2] & ~S[1] & ~S[0] & ~A[1] & ~A[0] //S4 -- 00
							| ~S[3] & S[2] & ~S[1] & S[0] & A[1] & A[0] //S5 -- 11
							| ~S[3] & S[2] & S[1] & S[0] & A[1] & ~A[0] //S7 -- 10
							| S[3] & ~S[2] & ~S[1] & ~S[0] & ~A[1] & A[0]; //S8 -- 01
							
	assign S_next[5] = ~S[3] & ~S[2] & ~S[1] & S[0] & A[1] & A[0] //S1 -- 11
							| ~S[3] & ~S[2] & S[1] & S[0] & A[1] & ~A[0] //S3 -- 10
							| ~S[3] & S[2] & ~S[1] & ~S[0] & ~A[1] & A[0] //S4 -- 01
							| ~S[3] & S[2] & S[1] & ~S[0] & A[1] & A[0] //S6 -- 11
							| S[3] & ~S[2] & ~S[1] & ~S[0] & A[1] & ~A[0]; //S8 -- 10
	
	assign S_next[6] = ~S[3] & ~S[2] & S[1] & ~S[0] & A[1] & A[0] //S2 -- 11
							| ~S[3] & S[2] & ~S[1] & ~S[0] & A[1] & ~A[0] //S4 -- 10
							| ~S[3] & S[2] & S[1] & S[0] & A[1] & A[0]; //S7 -- 11
	
	assign S_next[7] = ~S[3] & ~S[2] & S[1] & S[0] & A[1] & A[0] //S3 -- 11
							| S[3] & ~S[2] & ~S[1] & ~S[0] & A[1] & A[0]; //S8 -- 11
	
	assign S_next[8] = ~S[3] & S[2] & ~S[1] & ~S[0] & A[1] & A[0]; //S4 -- 11
	
	
	//Send the bits out based on state
	assign Out[0] = S_next[1] | S_next[3] | S_next[5] | S_next[7];
	assign Out[1] = S_next[2] | S_next[3] | S_next[6] | S_next[7];
	assign Out[2] = S_next[4] | S_next[5] | S_next[6] | S_next[7];
	assign Out[3] = S_next[8];
	
endmodule